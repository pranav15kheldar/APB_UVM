package apb_pkg;
 import uvm_pkg::*;
 `include "uvm_macros.svh"
 //`include "apb_interface.sv"
 `include "apb_seq_item.sv"
 `include "apb_seq_item_new.sv"
 `include "PrimeAddress_seq_item.sv"
 `include "apb_base_seq.sv" 
 `include "apb_seq.sv" 
 `include "apb_seq_read.sv"
 `include "PrimeAddress_sequence.sv" 
 `include "apb_sequencer.sv" 
 `include "apb_driver.sv" 
 `include "apb_agent.sv" 
 `include "apb_env.sv" 
 `include "apb_test.sv" 
 `include "PrimeAddress_test.sv"
endpackage
